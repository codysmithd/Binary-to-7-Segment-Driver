case "0000000000" => BCD_output <= "000000000000001111110";
case "0000000001" => BCD_output <= "000000000000000110000";
case "0000000010" => BCD_output <= "000000000000001101101";
case "0000000011" => BCD_output <= "000000000000001111001";
case "0000000100" => BCD_output <= "000000000000000110011";
case "0000000101" => BCD_output <= "000000000000001011011";
case "0000000110" => BCD_output <= "000000000000001011111";
case "0000000111" => BCD_output <= "000000000000001110000";
case "0000001000" => BCD_output <= "000000000000001111111";
case "0000001001" => BCD_output <= "000000000000001111011";
case "0000001010" => BCD_output <= "000000001100001111110";
case "0000001011" => BCD_output <= "000000001100000110000";
case "0000001100" => BCD_output <= "000000001100001101101";
case "0000001101" => BCD_output <= "000000001100001111001";
case "0000001110" => BCD_output <= "000000001100000110011";
case "0000001111" => BCD_output <= "000000001100001011011";
case "0000010000" => BCD_output <= "000000001100001011111";
case "0000010001" => BCD_output <= "000000001100001110000";
case "0000010010" => BCD_output <= "000000001100001111111";
case "0000010011" => BCD_output <= "000000001100001111011";
case "0000010100" => BCD_output <= "000000011011011111110";
case "0000010101" => BCD_output <= "000000011011010110000";
case "0000010110" => BCD_output <= "000000011011011101101";
case "0000010111" => BCD_output <= "000000011011011111001";
case "0000011000" => BCD_output <= "000000011011010110011";
case "0000011001" => BCD_output <= "000000011011011011011";
case "0000011010" => BCD_output <= "000000011011011011111";
case "0000011011" => BCD_output <= "000000011011011110000";
case "0000011100" => BCD_output <= "000000011011011111111";
case "0000011101" => BCD_output <= "000000011011011111011";
case "0000011110" => BCD_output <= "000000011110011111110";
case "0000011111" => BCD_output <= "000000011110010110000";
case "0000100000" => BCD_output <= "000000011110011101101";
case "0000100001" => BCD_output <= "000000011110011111001";
case "0000100010" => BCD_output <= "000000011110010110011";
case "0000100011" => BCD_output <= "000000011110011011011";
case "0000100100" => BCD_output <= "000000011110011011111";
case "0000100101" => BCD_output <= "000000011110011110000";
case "0000100110" => BCD_output <= "000000011110011111111";
case "0000100111" => BCD_output <= "000000011110011111011";
case "0000101000" => BCD_output <= "000000001100111111110";
case "0000101001" => BCD_output <= "000000001100110110000";
case "0000101010" => BCD_output <= "000000001100111101101";
case "0000101011" => BCD_output <= "000000001100111111001";
case "0000101100" => BCD_output <= "000000001100110110011";
case "0000101101" => BCD_output <= "000000001100111011011";
case "0000101110" => BCD_output <= "000000001100111011111";
case "0000101111" => BCD_output <= "000000001100111110000";
case "0000110000" => BCD_output <= "000000001100111111111";
case "0000110001" => BCD_output <= "000000001100111111011";
case "0000110010" => BCD_output <= "000000010110111111110";
case "0000110011" => BCD_output <= "000000010110110110000";
case "0000110100" => BCD_output <= "000000010110111101101";
case "0000110101" => BCD_output <= "000000010110111111001";
case "0000110110" => BCD_output <= "000000010110110110011";
case "0000110111" => BCD_output <= "000000010110111011011";
case "0000111000" => BCD_output <= "000000010110111011111";
case "0000111001" => BCD_output <= "000000010110111110000";
case "0000111010" => BCD_output <= "000000010110111111111";
case "0000111011" => BCD_output <= "000000010110111111011";
case "0000111100" => BCD_output <= "000000010111111111110";
case "0000111101" => BCD_output <= "000000010111110110000";
case "0000111110" => BCD_output <= "000000010111111101101";
case "0000111111" => BCD_output <= "000000010111111111001";
case "0001000000" => BCD_output <= "000000010111110110011";
case "0001000001" => BCD_output <= "000000010111111011011";
case "0001000010" => BCD_output <= "000000010111111011111";
case "0001000011" => BCD_output <= "000000010111111110000";
case "0001000100" => BCD_output <= "000000010111111111111";
case "0001000101" => BCD_output <= "000000010111111111011";
case "0001000110" => BCD_output <= "000000011100001111110";
case "0001000111" => BCD_output <= "000000011100000110000";
case "0001001000" => BCD_output <= "000000011100001101101";
case "0001001001" => BCD_output <= "000000011100001111001";
case "0001001010" => BCD_output <= "000000011100000110011";
case "0001001011" => BCD_output <= "000000011100001011011";
case "0001001100" => BCD_output <= "000000011100001011111";
case "0001001101" => BCD_output <= "000000011100001110000";
case "0001001110" => BCD_output <= "000000011100001111111";
case "0001001111" => BCD_output <= "000000011100001111011";
case "0001010000" => BCD_output <= "000000011111111111110";
case "0001010001" => BCD_output <= "000000011111110110000";
case "0001010010" => BCD_output <= "000000011111111101101";
case "0001010011" => BCD_output <= "000000011111111111001";
case "0001010100" => BCD_output <= "000000011111110110011";
case "0001010101" => BCD_output <= "000000011111111011011";
case "0001010110" => BCD_output <= "000000011111111011111";
case "0001010111" => BCD_output <= "000000011111111110000";
case "0001011000" => BCD_output <= "000000011111111111111";
case "0001011001" => BCD_output <= "000000011111111111011";
case "0001011010" => BCD_output <= "000000011110111111110";
case "0001011011" => BCD_output <= "000000011110110110000";
case "0001011100" => BCD_output <= "000000011110111101101";
case "0001011101" => BCD_output <= "000000011110111111001";
case "0001011110" => BCD_output <= "000000011110110110011";
case "0001011111" => BCD_output <= "000000011110111011011";
case "0001100000" => BCD_output <= "000000011110111011111";
case "0001100001" => BCD_output <= "000000011110111110000";
case "0001100010" => BCD_output <= "000000011110111111111";
case "0001100011" => BCD_output <= "000000011110111111011";
case "0001100100" => BCD_output <= "011000011111101111110";
case "0001100101" => BCD_output <= "011000011111100110000";
case "0001100110" => BCD_output <= "011000011111101101101";
case "0001100111" => BCD_output <= "011000011111101111001";
case "0001101000" => BCD_output <= "011000011111100110011";
case "0001101001" => BCD_output <= "011000011111101011011";
case "0001101010" => BCD_output <= "011000011111101011111";
case "0001101011" => BCD_output <= "011000011111101110000";
case "0001101100" => BCD_output <= "011000011111101111111";
case "0001101101" => BCD_output <= "011000011111101111011";
case "0001101110" => BCD_output <= "011000001100001111110";
case "0001101111" => BCD_output <= "011000001100000110000";
case "0001110000" => BCD_output <= "011000001100001101101";
case "0001110001" => BCD_output <= "011000001100001111001";
case "0001110010" => BCD_output <= "011000001100000110011";
case "0001110011" => BCD_output <= "011000001100001011011";
case "0001110100" => BCD_output <= "011000001100001011111";
case "0001110101" => BCD_output <= "011000001100001110000";
case "0001110110" => BCD_output <= "011000001100001111111";
case "0001110111" => BCD_output <= "011000001100001111011";
case "0001111000" => BCD_output <= "011000011011011111110";
case "0001111001" => BCD_output <= "011000011011010110000";
case "0001111010" => BCD_output <= "011000011011011101101";
case "0001111011" => BCD_output <= "011000011011011111001";
case "0001111100" => BCD_output <= "011000011011010110011";
case "0001111101" => BCD_output <= "011000011011011011011";
case "0001111110" => BCD_output <= "011000011011011011111";
case "0001111111" => BCD_output <= "011000011011011110000";
case "0010000000" => BCD_output <= "011000011011011111111";
case "0010000001" => BCD_output <= "011000011011011111011";
case "0010000010" => BCD_output <= "011000011110011111110";
case "0010000011" => BCD_output <= "011000011110010110000";
case "0010000100" => BCD_output <= "011000011110011101101";
case "0010000101" => BCD_output <= "011000011110011111001";
case "0010000110" => BCD_output <= "011000011110010110011";
case "0010000111" => BCD_output <= "011000011110011011011";
case "0010001000" => BCD_output <= "011000011110011011111";
case "0010001001" => BCD_output <= "011000011110011110000";
case "0010001010" => BCD_output <= "011000011110011111111";
case "0010001011" => BCD_output <= "011000011110011111011";
case "0010001100" => BCD_output <= "011000001100111111110";
case "0010001101" => BCD_output <= "011000001100110110000";
case "0010001110" => BCD_output <= "011000001100111101101";
case "0010001111" => BCD_output <= "011000001100111111001";
case "0010010000" => BCD_output <= "011000001100110110011";
case "0010010001" => BCD_output <= "011000001100111011011";
case "0010010010" => BCD_output <= "011000001100111011111";
case "0010010011" => BCD_output <= "011000001100111110000";
case "0010010100" => BCD_output <= "011000001100111111111";
case "0010010101" => BCD_output <= "011000001100111111011";
case "0010010110" => BCD_output <= "011000010110111111110";
case "0010010111" => BCD_output <= "011000010110110110000";
case "0010011000" => BCD_output <= "011000010110111101101";
case "0010011001" => BCD_output <= "011000010110111111001";
case "0010011010" => BCD_output <= "011000010110110110011";
case "0010011011" => BCD_output <= "011000010110111011011";
case "0010011100" => BCD_output <= "011000010110111011111";
case "0010011101" => BCD_output <= "011000010110111110000";
case "0010011110" => BCD_output <= "011000010110111111111";
case "0010011111" => BCD_output <= "011000010110111111011";
case "0010100000" => BCD_output <= "011000010111111111110";
case "0010100001" => BCD_output <= "011000010111110110000";
case "0010100010" => BCD_output <= "011000010111111101101";
case "0010100011" => BCD_output <= "011000010111111111001";
case "0010100100" => BCD_output <= "011000010111110110011";
case "0010100101" => BCD_output <= "011000010111111011011";
case "0010100110" => BCD_output <= "011000010111111011111";
case "0010100111" => BCD_output <= "011000010111111110000";
case "0010101000" => BCD_output <= "011000010111111111111";
case "0010101001" => BCD_output <= "011000010111111111011";
case "0010101010" => BCD_output <= "011000011100001111110";
case "0010101011" => BCD_output <= "011000011100000110000";
case "0010101100" => BCD_output <= "011000011100001101101";
case "0010101101" => BCD_output <= "011000011100001111001";
case "0010101110" => BCD_output <= "011000011100000110011";
case "0010101111" => BCD_output <= "011000011100001011011";
case "0010110000" => BCD_output <= "011000011100001011111";
case "0010110001" => BCD_output <= "011000011100001110000";
case "0010110010" => BCD_output <= "011000011100001111111";
case "0010110011" => BCD_output <= "011000011100001111011";
case "0010110100" => BCD_output <= "011000011111111111110";
case "0010110101" => BCD_output <= "011000011111110110000";
case "0010110110" => BCD_output <= "011000011111111101101";
case "0010110111" => BCD_output <= "011000011111111111001";
case "0010111000" => BCD_output <= "011000011111110110011";
case "0010111001" => BCD_output <= "011000011111111011011";
case "0010111010" => BCD_output <= "011000011111111011111";
case "0010111011" => BCD_output <= "011000011111111110000";
case "0010111100" => BCD_output <= "011000011111111111111";
case "0010111101" => BCD_output <= "011000011111111111011";
case "0010111110" => BCD_output <= "011000011110111111110";
case "0010111111" => BCD_output <= "011000011110110110000";
case "0011000000" => BCD_output <= "011000011110111101101";
case "0011000001" => BCD_output <= "011000011110111111001";
case "0011000010" => BCD_output <= "011000011110110110011";
case "0011000011" => BCD_output <= "011000011110111011011";
case "0011000100" => BCD_output <= "011000011110111011111";
case "0011000101" => BCD_output <= "011000011110111110000";
case "0011000110" => BCD_output <= "011000011110111111111";
case "0011000111" => BCD_output <= "011000011110111111011";
case "0011001000" => BCD_output <= "110110111111101111110";
case "0011001001" => BCD_output <= "110110111111100110000";
case "0011001010" => BCD_output <= "110110111111101101101";
case "0011001011" => BCD_output <= "110110111111101111001";
case "0011001100" => BCD_output <= "110110111111100110011";
case "0011001101" => BCD_output <= "110110111111101011011";
case "0011001110" => BCD_output <= "110110111111101011111";
case "0011001111" => BCD_output <= "110110111111101110000";
case "0011010000" => BCD_output <= "110110111111101111111";
case "0011010001" => BCD_output <= "110110111111101111011";
case "0011010010" => BCD_output <= "110110101100001111110";
case "0011010011" => BCD_output <= "110110101100000110000";
case "0011010100" => BCD_output <= "110110101100001101101";
case "0011010101" => BCD_output <= "110110101100001111001";
case "0011010110" => BCD_output <= "110110101100000110011";
case "0011010111" => BCD_output <= "110110101100001011011";
case "0011011000" => BCD_output <= "110110101100001011111";
case "0011011001" => BCD_output <= "110110101100001110000";
case "0011011010" => BCD_output <= "110110101100001111111";
case "0011011011" => BCD_output <= "110110101100001111011";
case "0011011100" => BCD_output <= "110110111011011111110";
case "0011011101" => BCD_output <= "110110111011010110000";
case "0011011110" => BCD_output <= "110110111011011101101";
case "0011011111" => BCD_output <= "110110111011011111001";
case "0011100000" => BCD_output <= "110110111011010110011";
case "0011100001" => BCD_output <= "110110111011011011011";
case "0011100010" => BCD_output <= "110110111011011011111";
case "0011100011" => BCD_output <= "110110111011011110000";
case "0011100100" => BCD_output <= "110110111011011111111";
case "0011100101" => BCD_output <= "110110111011011111011";
case "0011100110" => BCD_output <= "110110111110011111110";
case "0011100111" => BCD_output <= "110110111110010110000";
case "0011101000" => BCD_output <= "110110111110011101101";
case "0011101001" => BCD_output <= "110110111110011111001";
case "0011101010" => BCD_output <= "110110111110010110011";
case "0011101011" => BCD_output <= "110110111110011011011";
case "0011101100" => BCD_output <= "110110111110011011111";
case "0011101101" => BCD_output <= "110110111110011110000";
case "0011101110" => BCD_output <= "110110111110011111111";
case "0011101111" => BCD_output <= "110110111110011111011";
case "0011110000" => BCD_output <= "110110101100111111110";
case "0011110001" => BCD_output <= "110110101100110110000";
case "0011110010" => BCD_output <= "110110101100111101101";
case "0011110011" => BCD_output <= "110110101100111111001";
case "0011110100" => BCD_output <= "110110101100110110011";
case "0011110101" => BCD_output <= "110110101100111011011";
case "0011110110" => BCD_output <= "110110101100111011111";
case "0011110111" => BCD_output <= "110110101100111110000";
case "0011111000" => BCD_output <= "110110101100111111111";
case "0011111001" => BCD_output <= "110110101100111111011";
case "0011111010" => BCD_output <= "110110110110111111110";
case "0011111011" => BCD_output <= "110110110110110110000";
case "0011111100" => BCD_output <= "110110110110111101101";
case "0011111101" => BCD_output <= "110110110110111111001";
case "0011111110" => BCD_output <= "110110110110110110011";
case "0011111111" => BCD_output <= "110110110110111011011";
case "0100000000" => BCD_output <= "110110110110111011111";
case "0100000001" => BCD_output <= "110110110110111110000";
case "0100000010" => BCD_output <= "110110110110111111111";
case "0100000011" => BCD_output <= "110110110110111111011";
case "0100000100" => BCD_output <= "110110110111111111110";
case "0100000101" => BCD_output <= "110110110111110110000";
case "0100000110" => BCD_output <= "110110110111111101101";
case "0100000111" => BCD_output <= "110110110111111111001";
case "0100001000" => BCD_output <= "110110110111110110011";
case "0100001001" => BCD_output <= "110110110111111011011";
case "0100001010" => BCD_output <= "110110110111111011111";
case "0100001011" => BCD_output <= "110110110111111110000";
case "0100001100" => BCD_output <= "110110110111111111111";
case "0100001101" => BCD_output <= "110110110111111111011";
case "0100001110" => BCD_output <= "110110111100001111110";
case "0100001111" => BCD_output <= "110110111100000110000";
case "0100010000" => BCD_output <= "110110111100001101101";
case "0100010001" => BCD_output <= "110110111100001111001";
case "0100010010" => BCD_output <= "110110111100000110011";
case "0100010011" => BCD_output <= "110110111100001011011";
case "0100010100" => BCD_output <= "110110111100001011111";
case "0100010101" => BCD_output <= "110110111100001110000";
case "0100010110" => BCD_output <= "110110111100001111111";
case "0100010111" => BCD_output <= "110110111100001111011";
case "0100011000" => BCD_output <= "110110111111111111110";
case "0100011001" => BCD_output <= "110110111111110110000";
case "0100011010" => BCD_output <= "110110111111111101101";
case "0100011011" => BCD_output <= "110110111111111111001";
case "0100011100" => BCD_output <= "110110111111110110011";
case "0100011101" => BCD_output <= "110110111111111011011";
case "0100011110" => BCD_output <= "110110111111111011111";
case "0100011111" => BCD_output <= "110110111111111110000";
case "0100100000" => BCD_output <= "110110111111111111111";
case "0100100001" => BCD_output <= "110110111111111111011";
case "0100100010" => BCD_output <= "110110111110111111110";
case "0100100011" => BCD_output <= "110110111110110110000";
case "0100100100" => BCD_output <= "110110111110111101101";
case "0100100101" => BCD_output <= "110110111110111111001";
case "0100100110" => BCD_output <= "110110111110110110011";
case "0100100111" => BCD_output <= "110110111110111011011";
case "0100101000" => BCD_output <= "110110111110111011111";
case "0100101001" => BCD_output <= "110110111110111110000";
case "0100101010" => BCD_output <= "110110111110111111111";
case "0100101011" => BCD_output <= "110110111110111111011";
case "0100101100" => BCD_output <= "111100111111101111110";
case "0100101101" => BCD_output <= "111100111111100110000";
case "0100101110" => BCD_output <= "111100111111101101101";
case "0100101111" => BCD_output <= "111100111111101111001";
case "0100110000" => BCD_output <= "111100111111100110011";
case "0100110001" => BCD_output <= "111100111111101011011";
case "0100110010" => BCD_output <= "111100111111101011111";
case "0100110011" => BCD_output <= "111100111111101110000";
case "0100110100" => BCD_output <= "111100111111101111111";
case "0100110101" => BCD_output <= "111100111111101111011";
case "0100110110" => BCD_output <= "111100101100001111110";
case "0100110111" => BCD_output <= "111100101100000110000";
case "0100111000" => BCD_output <= "111100101100001101101";
case "0100111001" => BCD_output <= "111100101100001111001";
case "0100111010" => BCD_output <= "111100101100000110011";
case "0100111011" => BCD_output <= "111100101100001011011";
case "0100111100" => BCD_output <= "111100101100001011111";
case "0100111101" => BCD_output <= "111100101100001110000";
case "0100111110" => BCD_output <= "111100101100001111111";
case "0100111111" => BCD_output <= "111100101100001111011";
case "0101000000" => BCD_output <= "111100111011011111110";
case "0101000001" => BCD_output <= "111100111011010110000";
case "0101000010" => BCD_output <= "111100111011011101101";
case "0101000011" => BCD_output <= "111100111011011111001";
case "0101000100" => BCD_output <= "111100111011010110011";
case "0101000101" => BCD_output <= "111100111011011011011";
case "0101000110" => BCD_output <= "111100111011011011111";
case "0101000111" => BCD_output <= "111100111011011110000";
case "0101001000" => BCD_output <= "111100111011011111111";
case "0101001001" => BCD_output <= "111100111011011111011";
case "0101001010" => BCD_output <= "111100111110011111110";
case "0101001011" => BCD_output <= "111100111110010110000";
case "0101001100" => BCD_output <= "111100111110011101101";
case "0101001101" => BCD_output <= "111100111110011111001";
case "0101001110" => BCD_output <= "111100111110010110011";
case "0101001111" => BCD_output <= "111100111110011011011";
case "0101010000" => BCD_output <= "111100111110011011111";
case "0101010001" => BCD_output <= "111100111110011110000";
case "0101010010" => BCD_output <= "111100111110011111111";
case "0101010011" => BCD_output <= "111100111110011111011";
case "0101010100" => BCD_output <= "111100101100111111110";
case "0101010101" => BCD_output <= "111100101100110110000";
case "0101010110" => BCD_output <= "111100101100111101101";
case "0101010111" => BCD_output <= "111100101100111111001";
case "0101011000" => BCD_output <= "111100101100110110011";
case "0101011001" => BCD_output <= "111100101100111011011";
case "0101011010" => BCD_output <= "111100101100111011111";
case "0101011011" => BCD_output <= "111100101100111110000";
case "0101011100" => BCD_output <= "111100101100111111111";
case "0101011101" => BCD_output <= "111100101100111111011";
case "0101011110" => BCD_output <= "111100110110111111110";
case "0101011111" => BCD_output <= "111100110110110110000";
case "0101100000" => BCD_output <= "111100110110111101101";
case "0101100001" => BCD_output <= "111100110110111111001";
case "0101100010" => BCD_output <= "111100110110110110011";
case "0101100011" => BCD_output <= "111100110110111011011";
case "0101100100" => BCD_output <= "111100110110111011111";
case "0101100101" => BCD_output <= "111100110110111110000";
case "0101100110" => BCD_output <= "111100110110111111111";
case "0101100111" => BCD_output <= "111100110110111111011";
case "0101101000" => BCD_output <= "111100110111111111110";
case "0101101001" => BCD_output <= "111100110111110110000";
case "0101101010" => BCD_output <= "111100110111111101101";
case "0101101011" => BCD_output <= "111100110111111111001";
case "0101101100" => BCD_output <= "111100110111110110011";
case "0101101101" => BCD_output <= "111100110111111011011";
case "0101101110" => BCD_output <= "111100110111111011111";
case "0101101111" => BCD_output <= "111100110111111110000";
case "0101110000" => BCD_output <= "111100110111111111111";
case "0101110001" => BCD_output <= "111100110111111111011";
case "0101110010" => BCD_output <= "111100111100001111110";
case "0101110011" => BCD_output <= "111100111100000110000";
case "0101110100" => BCD_output <= "111100111100001101101";
case "0101110101" => BCD_output <= "111100111100001111001";
case "0101110110" => BCD_output <= "111100111100000110011";
case "0101110111" => BCD_output <= "111100111100001011011";
case "0101111000" => BCD_output <= "111100111100001011111";
case "0101111001" => BCD_output <= "111100111100001110000";
case "0101111010" => BCD_output <= "111100111100001111111";
case "0101111011" => BCD_output <= "111100111100001111011";
case "0101111100" => BCD_output <= "111100111111111111110";
case "0101111101" => BCD_output <= "111100111111110110000";
case "0101111110" => BCD_output <= "111100111111111101101";
case "0101111111" => BCD_output <= "111100111111111111001";
case "0110000000" => BCD_output <= "111100111111110110011";
case "0110000001" => BCD_output <= "111100111111111011011";
case "0110000010" => BCD_output <= "111100111111111011111";
case "0110000011" => BCD_output <= "111100111111111110000";
case "0110000100" => BCD_output <= "111100111111111111111";
case "0110000101" => BCD_output <= "111100111111111111011";
case "0110000110" => BCD_output <= "111100111110111111110";
case "0110000111" => BCD_output <= "111100111110110110000";
case "0110001000" => BCD_output <= "111100111110111101101";
case "0110001001" => BCD_output <= "111100111110111111001";
case "0110001010" => BCD_output <= "111100111110110110011";
case "0110001011" => BCD_output <= "111100111110111011011";
case "0110001100" => BCD_output <= "111100111110111011111";
case "0110001101" => BCD_output <= "111100111110111110000";
case "0110001110" => BCD_output <= "111100111110111111111";
case "0110001111" => BCD_output <= "111100111110111111011";
case "0110010000" => BCD_output <= "011001111111101111110";
case "0110010001" => BCD_output <= "011001111111100110000";
case "0110010010" => BCD_output <= "011001111111101101101";
case "0110010011" => BCD_output <= "011001111111101111001";
case "0110010100" => BCD_output <= "011001111111100110011";
case "0110010101" => BCD_output <= "011001111111101011011";
case "0110010110" => BCD_output <= "011001111111101011111";
case "0110010111" => BCD_output <= "011001111111101110000";
case "0110011000" => BCD_output <= "011001111111101111111";
case "0110011001" => BCD_output <= "011001111111101111011";
case "0110011010" => BCD_output <= "011001101100001111110";
case "0110011011" => BCD_output <= "011001101100000110000";
case "0110011100" => BCD_output <= "011001101100001101101";
case "0110011101" => BCD_output <= "011001101100001111001";
case "0110011110" => BCD_output <= "011001101100000110011";
case "0110011111" => BCD_output <= "011001101100001011011";
case "0110100000" => BCD_output <= "011001101100001011111";
case "0110100001" => BCD_output <= "011001101100001110000";
case "0110100010" => BCD_output <= "011001101100001111111";
case "0110100011" => BCD_output <= "011001101100001111011";
case "0110100100" => BCD_output <= "011001111011011111110";
case "0110100101" => BCD_output <= "011001111011010110000";
case "0110100110" => BCD_output <= "011001111011011101101";
case "0110100111" => BCD_output <= "011001111011011111001";
case "0110101000" => BCD_output <= "011001111011010110011";
case "0110101001" => BCD_output <= "011001111011011011011";
case "0110101010" => BCD_output <= "011001111011011011111";
case "0110101011" => BCD_output <= "011001111011011110000";
case "0110101100" => BCD_output <= "011001111011011111111";
case "0110101101" => BCD_output <= "011001111011011111011";
case "0110101110" => BCD_output <= "011001111110011111110";
case "0110101111" => BCD_output <= "011001111110010110000";
case "0110110000" => BCD_output <= "011001111110011101101";
case "0110110001" => BCD_output <= "011001111110011111001";
case "0110110010" => BCD_output <= "011001111110010110011";
case "0110110011" => BCD_output <= "011001111110011011011";
case "0110110100" => BCD_output <= "011001111110011011111";
case "0110110101" => BCD_output <= "011001111110011110000";
case "0110110110" => BCD_output <= "011001111110011111111";
case "0110110111" => BCD_output <= "011001111110011111011";
case "0110111000" => BCD_output <= "011001101100111111110";
case "0110111001" => BCD_output <= "011001101100110110000";
case "0110111010" => BCD_output <= "011001101100111101101";
case "0110111011" => BCD_output <= "011001101100111111001";
case "0110111100" => BCD_output <= "011001101100110110011";
case "0110111101" => BCD_output <= "011001101100111011011";
case "0110111110" => BCD_output <= "011001101100111011111";
case "0110111111" => BCD_output <= "011001101100111110000";
case "0111000000" => BCD_output <= "011001101100111111111";
case "0111000001" => BCD_output <= "011001101100111111011";
case "0111000010" => BCD_output <= "011001110110111111110";
case "0111000011" => BCD_output <= "011001110110110110000";
case "0111000100" => BCD_output <= "011001110110111101101";
case "0111000101" => BCD_output <= "011001110110111111001";
case "0111000110" => BCD_output <= "011001110110110110011";
case "0111000111" => BCD_output <= "011001110110111011011";
case "0111001000" => BCD_output <= "011001110110111011111";
case "0111001001" => BCD_output <= "011001110110111110000";
case "0111001010" => BCD_output <= "011001110110111111111";
case "0111001011" => BCD_output <= "011001110110111111011";
case "0111001100" => BCD_output <= "011001110111111111110";
case "0111001101" => BCD_output <= "011001110111110110000";
case "0111001110" => BCD_output <= "011001110111111101101";
case "0111001111" => BCD_output <= "011001110111111111001";
case "0111010000" => BCD_output <= "011001110111110110011";
case "0111010001" => BCD_output <= "011001110111111011011";
case "0111010010" => BCD_output <= "011001110111111011111";
case "0111010011" => BCD_output <= "011001110111111110000";
case "0111010100" => BCD_output <= "011001110111111111111";
case "0111010101" => BCD_output <= "011001110111111111011";
case "0111010110" => BCD_output <= "011001111100001111110";
case "0111010111" => BCD_output <= "011001111100000110000";
case "0111011000" => BCD_output <= "011001111100001101101";
case "0111011001" => BCD_output <= "011001111100001111001";
case "0111011010" => BCD_output <= "011001111100000110011";
case "0111011011" => BCD_output <= "011001111100001011011";
case "0111011100" => BCD_output <= "011001111100001011111";
case "0111011101" => BCD_output <= "011001111100001110000";
case "0111011110" => BCD_output <= "011001111100001111111";
case "0111011111" => BCD_output <= "011001111100001111011";
case "0111100000" => BCD_output <= "011001111111111111110";
case "0111100001" => BCD_output <= "011001111111110110000";
case "0111100010" => BCD_output <= "011001111111111101101";
case "0111100011" => BCD_output <= "011001111111111111001";
case "0111100100" => BCD_output <= "011001111111110110011";
case "0111100101" => BCD_output <= "011001111111111011011";
case "0111100110" => BCD_output <= "011001111111111011111";
case "0111100111" => BCD_output <= "011001111111111110000";
case "0111101000" => BCD_output <= "011001111111111111111";
case "0111101001" => BCD_output <= "011001111111111111011";
case "0111101010" => BCD_output <= "011001111110111111110";
case "0111101011" => BCD_output <= "011001111110110110000";
case "0111101100" => BCD_output <= "011001111110111101101";
case "0111101101" => BCD_output <= "011001111110111111001";
case "0111101110" => BCD_output <= "011001111110110110011";
case "0111101111" => BCD_output <= "011001111110111011011";
case "0111110000" => BCD_output <= "011001111110111011111";
case "0111110001" => BCD_output <= "011001111110111110000";
case "0111110010" => BCD_output <= "011001111110111111111";
case "0111110011" => BCD_output <= "011001111110111111011";
case "0111110100" => BCD_output <= "101101111111101111110";
case "0111110101" => BCD_output <= "101101111111100110000";
case "0111110110" => BCD_output <= "101101111111101101101";
case "0111110111" => BCD_output <= "101101111111101111001";
case "0111111000" => BCD_output <= "101101111111100110011";
case "0111111001" => BCD_output <= "101101111111101011011";
case "0111111010" => BCD_output <= "101101111111101011111";
case "0111111011" => BCD_output <= "101101111111101110000";
case "0111111100" => BCD_output <= "101101111111101111111";
case "0111111101" => BCD_output <= "101101111111101111011";
case "0111111110" => BCD_output <= "101101101100001111110";
case "0111111111" => BCD_output <= "101101101100000110000";
case "1000000000" => BCD_output <= "101101101100001101101";
case "1000000001" => BCD_output <= "101101101100001111001";
case "1000000010" => BCD_output <= "101101101100000110011";
case "1000000011" => BCD_output <= "101101101100001011011";
case "1000000100" => BCD_output <= "101101101100001011111";
case "1000000101" => BCD_output <= "101101101100001110000";
case "1000000110" => BCD_output <= "101101101100001111111";
case "1000000111" => BCD_output <= "101101101100001111011";
case "1000001000" => BCD_output <= "101101111011011111110";
case "1000001001" => BCD_output <= "101101111011010110000";
case "1000001010" => BCD_output <= "101101111011011101101";
case "1000001011" => BCD_output <= "101101111011011111001";
case "1000001100" => BCD_output <= "101101111011010110011";
case "1000001101" => BCD_output <= "101101111011011011011";
case "1000001110" => BCD_output <= "101101111011011011111";
case "1000001111" => BCD_output <= "101101111011011110000";
case "1000010000" => BCD_output <= "101101111011011111111";
case "1000010001" => BCD_output <= "101101111011011111011";
case "1000010010" => BCD_output <= "101101111110011111110";
case "1000010011" => BCD_output <= "101101111110010110000";
case "1000010100" => BCD_output <= "101101111110011101101";
case "1000010101" => BCD_output <= "101101111110011111001";
case "1000010110" => BCD_output <= "101101111110010110011";
case "1000010111" => BCD_output <= "101101111110011011011";
case "1000011000" => BCD_output <= "101101111110011011111";
case "1000011001" => BCD_output <= "101101111110011110000";
case "1000011010" => BCD_output <= "101101111110011111111";
case "1000011011" => BCD_output <= "101101111110011111011";
case "1000011100" => BCD_output <= "101101101100111111110";
case "1000011101" => BCD_output <= "101101101100110110000";
case "1000011110" => BCD_output <= "101101101100111101101";
case "1000011111" => BCD_output <= "101101101100111111001";
case "1000100000" => BCD_output <= "101101101100110110011";
case "1000100001" => BCD_output <= "101101101100111011011";
case "1000100010" => BCD_output <= "101101101100111011111";
case "1000100011" => BCD_output <= "101101101100111110000";
case "1000100100" => BCD_output <= "101101101100111111111";
case "1000100101" => BCD_output <= "101101101100111111011";
case "1000100110" => BCD_output <= "101101110110111111110";
case "1000100111" => BCD_output <= "101101110110110110000";
case "1000101000" => BCD_output <= "101101110110111101101";
case "1000101001" => BCD_output <= "101101110110111111001";
case "1000101010" => BCD_output <= "101101110110110110011";
case "1000101011" => BCD_output <= "101101110110111011011";
case "1000101100" => BCD_output <= "101101110110111011111";
case "1000101101" => BCD_output <= "101101110110111110000";
case "1000101110" => BCD_output <= "101101110110111111111";
case "1000101111" => BCD_output <= "101101110110111111011";
case "1000110000" => BCD_output <= "101101110111111111110";
case "1000110001" => BCD_output <= "101101110111110110000";
case "1000110010" => BCD_output <= "101101110111111101101";
case "1000110011" => BCD_output <= "101101110111111111001";
case "1000110100" => BCD_output <= "101101110111110110011";
case "1000110101" => BCD_output <= "101101110111111011011";
case "1000110110" => BCD_output <= "101101110111111011111";
case "1000110111" => BCD_output <= "101101110111111110000";
case "1000111000" => BCD_output <= "101101110111111111111";
case "1000111001" => BCD_output <= "101101110111111111011";
case "1000111010" => BCD_output <= "101101111100001111110";
case "1000111011" => BCD_output <= "101101111100000110000";
case "1000111100" => BCD_output <= "101101111100001101101";
case "1000111101" => BCD_output <= "101101111100001111001";
case "1000111110" => BCD_output <= "101101111100000110011";
case "1000111111" => BCD_output <= "101101111100001011011";
case "1001000000" => BCD_output <= "101101111100001011111";
case "1001000001" => BCD_output <= "101101111100001110000";
case "1001000010" => BCD_output <= "101101111100001111111";
case "1001000011" => BCD_output <= "101101111100001111011";
case "1001000100" => BCD_output <= "101101111111111111110";
case "1001000101" => BCD_output <= "101101111111110110000";
case "1001000110" => BCD_output <= "101101111111111101101";
case "1001000111" => BCD_output <= "101101111111111111001";
case "1001001000" => BCD_output <= "101101111111110110011";
case "1001001001" => BCD_output <= "101101111111111011011";
case "1001001010" => BCD_output <= "101101111111111011111";
case "1001001011" => BCD_output <= "101101111111111110000";
case "1001001100" => BCD_output <= "101101111111111111111";
case "1001001101" => BCD_output <= "101101111111111111011";
case "1001001110" => BCD_output <= "101101111110111111110";
case "1001001111" => BCD_output <= "101101111110110110000";
case "1001010000" => BCD_output <= "101101111110111101101";
case "1001010001" => BCD_output <= "101101111110111111001";
case "1001010010" => BCD_output <= "101101111110110110011";
case "1001010011" => BCD_output <= "101101111110111011011";
case "1001010100" => BCD_output <= "101101111110111011111";
case "1001010101" => BCD_output <= "101101111110111110000";
case "1001010110" => BCD_output <= "101101111110111111111";
case "1001010111" => BCD_output <= "101101111110111111011";
case "1001011000" => BCD_output <= "101111111111101111110";
case "1001011001" => BCD_output <= "101111111111100110000";
case "1001011010" => BCD_output <= "101111111111101101101";
case "1001011011" => BCD_output <= "101111111111101111001";
case "1001011100" => BCD_output <= "101111111111100110011";
case "1001011101" => BCD_output <= "101111111111101011011";
case "1001011110" => BCD_output <= "101111111111101011111";
case "1001011111" => BCD_output <= "101111111111101110000";
case "1001100000" => BCD_output <= "101111111111101111111";
case "1001100001" => BCD_output <= "101111111111101111011";
case "1001100010" => BCD_output <= "101111101100001111110";
case "1001100011" => BCD_output <= "101111101100000110000";
case "1001100100" => BCD_output <= "101111101100001101101";
case "1001100101" => BCD_output <= "101111101100001111001";
case "1001100110" => BCD_output <= "101111101100000110011";
case "1001100111" => BCD_output <= "101111101100001011011";
case "1001101000" => BCD_output <= "101111101100001011111";
case "1001101001" => BCD_output <= "101111101100001110000";
case "1001101010" => BCD_output <= "101111101100001111111";
case "1001101011" => BCD_output <= "101111101100001111011";
case "1001101100" => BCD_output <= "101111111011011111110";
case "1001101101" => BCD_output <= "101111111011010110000";
case "1001101110" => BCD_output <= "101111111011011101101";
case "1001101111" => BCD_output <= "101111111011011111001";
case "1001110000" => BCD_output <= "101111111011010110011";
case "1001110001" => BCD_output <= "101111111011011011011";
case "1001110010" => BCD_output <= "101111111011011011111";
case "1001110011" => BCD_output <= "101111111011011110000";
case "1001110100" => BCD_output <= "101111111011011111111";
case "1001110101" => BCD_output <= "101111111011011111011";
case "1001110110" => BCD_output <= "101111111110011111110";
case "1001110111" => BCD_output <= "101111111110010110000";
case "1001111000" => BCD_output <= "101111111110011101101";
case "1001111001" => BCD_output <= "101111111110011111001";
case "1001111010" => BCD_output <= "101111111110010110011";
case "1001111011" => BCD_output <= "101111111110011011011";
case "1001111100" => BCD_output <= "101111111110011011111";
case "1001111101" => BCD_output <= "101111111110011110000";
case "1001111110" => BCD_output <= "101111111110011111111";
case "1001111111" => BCD_output <= "101111111110011111011";
case "1010000000" => BCD_output <= "101111101100111111110";
case "1010000001" => BCD_output <= "101111101100110110000";
case "1010000010" => BCD_output <= "101111101100111101101";
case "1010000011" => BCD_output <= "101111101100111111001";
case "1010000100" => BCD_output <= "101111101100110110011";
case "1010000101" => BCD_output <= "101111101100111011011";
case "1010000110" => BCD_output <= "101111101100111011111";
case "1010000111" => BCD_output <= "101111101100111110000";
case "1010001000" => BCD_output <= "101111101100111111111";
case "1010001001" => BCD_output <= "101111101100111111011";
case "1010001010" => BCD_output <= "101111110110111111110";
case "1010001011" => BCD_output <= "101111110110110110000";
case "1010001100" => BCD_output <= "101111110110111101101";
case "1010001101" => BCD_output <= "101111110110111111001";
case "1010001110" => BCD_output <= "101111110110110110011";
case "1010001111" => BCD_output <= "101111110110111011011";
case "1010010000" => BCD_output <= "101111110110111011111";
case "1010010001" => BCD_output <= "101111110110111110000";
case "1010010010" => BCD_output <= "101111110110111111111";
case "1010010011" => BCD_output <= "101111110110111111011";
case "1010010100" => BCD_output <= "101111110111111111110";
case "1010010101" => BCD_output <= "101111110111110110000";
case "1010010110" => BCD_output <= "101111110111111101101";
case "1010010111" => BCD_output <= "101111110111111111001";
case "1010011000" => BCD_output <= "101111110111110110011";
case "1010011001" => BCD_output <= "101111110111111011011";
case "1010011010" => BCD_output <= "101111110111111011111";
case "1010011011" => BCD_output <= "101111110111111110000";
case "1010011100" => BCD_output <= "101111110111111111111";
case "1010011101" => BCD_output <= "101111110111111111011";
case "1010011110" => BCD_output <= "101111111100001111110";
case "1010011111" => BCD_output <= "101111111100000110000";
case "1010100000" => BCD_output <= "101111111100001101101";
case "1010100001" => BCD_output <= "101111111100001111001";
case "1010100010" => BCD_output <= "101111111100000110011";
case "1010100011" => BCD_output <= "101111111100001011011";
case "1010100100" => BCD_output <= "101111111100001011111";
case "1010100101" => BCD_output <= "101111111100001110000";
case "1010100110" => BCD_output <= "101111111100001111111";
case "1010100111" => BCD_output <= "101111111100001111011";
case "1010101000" => BCD_output <= "101111111111111111110";
case "1010101001" => BCD_output <= "101111111111110110000";
case "1010101010" => BCD_output <= "101111111111111101101";
case "1010101011" => BCD_output <= "101111111111111111001";
case "1010101100" => BCD_output <= "101111111111110110011";
case "1010101101" => BCD_output <= "101111111111111011011";
case "1010101110" => BCD_output <= "101111111111111011111";
case "1010101111" => BCD_output <= "101111111111111110000";
case "1010110000" => BCD_output <= "101111111111111111111";
case "1010110001" => BCD_output <= "101111111111111111011";
case "1010110010" => BCD_output <= "101111111110111111110";
case "1010110011" => BCD_output <= "101111111110110110000";
case "1010110100" => BCD_output <= "101111111110111101101";
case "1010110101" => BCD_output <= "101111111110111111001";
case "1010110110" => BCD_output <= "101111111110110110011";
case "1010110111" => BCD_output <= "101111111110111011011";
case "1010111000" => BCD_output <= "101111111110111011111";
case "1010111001" => BCD_output <= "101111111110111110000";
case "1010111010" => BCD_output <= "101111111110111111111";
case "1010111011" => BCD_output <= "101111111110111111011";
case "1010111100" => BCD_output <= "111000011111101111110";
case "1010111101" => BCD_output <= "111000011111100110000";
case "1010111110" => BCD_output <= "111000011111101101101";
case "1010111111" => BCD_output <= "111000011111101111001";
case "1011000000" => BCD_output <= "111000011111100110011";
case "1011000001" => BCD_output <= "111000011111101011011";
case "1011000010" => BCD_output <= "111000011111101011111";
case "1011000011" => BCD_output <= "111000011111101110000";
case "1011000100" => BCD_output <= "111000011111101111111";
case "1011000101" => BCD_output <= "111000011111101111011";
case "1011000110" => BCD_output <= "111000001100001111110";
case "1011000111" => BCD_output <= "111000001100000110000";
case "1011001000" => BCD_output <= "111000001100001101101";
case "1011001001" => BCD_output <= "111000001100001111001";
case "1011001010" => BCD_output <= "111000001100000110011";
case "1011001011" => BCD_output <= "111000001100001011011";
case "1011001100" => BCD_output <= "111000001100001011111";
case "1011001101" => BCD_output <= "111000001100001110000";
case "1011001110" => BCD_output <= "111000001100001111111";
case "1011001111" => BCD_output <= "111000001100001111011";
case "1011010000" => BCD_output <= "111000011011011111110";
case "1011010001" => BCD_output <= "111000011011010110000";
case "1011010010" => BCD_output <= "111000011011011101101";
case "1011010011" => BCD_output <= "111000011011011111001";
case "1011010100" => BCD_output <= "111000011011010110011";
case "1011010101" => BCD_output <= "111000011011011011011";
case "1011010110" => BCD_output <= "111000011011011011111";
case "1011010111" => BCD_output <= "111000011011011110000";
case "1011011000" => BCD_output <= "111000011011011111111";
case "1011011001" => BCD_output <= "111000011011011111011";
case "1011011010" => BCD_output <= "111000011110011111110";
case "1011011011" => BCD_output <= "111000011110010110000";
case "1011011100" => BCD_output <= "111000011110011101101";
case "1011011101" => BCD_output <= "111000011110011111001";
case "1011011110" => BCD_output <= "111000011110010110011";
case "1011011111" => BCD_output <= "111000011110011011011";
case "1011100000" => BCD_output <= "111000011110011011111";
case "1011100001" => BCD_output <= "111000011110011110000";
case "1011100010" => BCD_output <= "111000011110011111111";
case "1011100011" => BCD_output <= "111000011110011111011";
case "1011100100" => BCD_output <= "111000001100111111110";
case "1011100101" => BCD_output <= "111000001100110110000";
case "1011100110" => BCD_output <= "111000001100111101101";
case "1011100111" => BCD_output <= "111000001100111111001";
case "1011101000" => BCD_output <= "111000001100110110011";
case "1011101001" => BCD_output <= "111000001100111011011";
case "1011101010" => BCD_output <= "111000001100111011111";
case "1011101011" => BCD_output <= "111000001100111110000";
case "1011101100" => BCD_output <= "111000001100111111111";
case "1011101101" => BCD_output <= "111000001100111111011";
case "1011101110" => BCD_output <= "111000010110111111110";
case "1011101111" => BCD_output <= "111000010110110110000";
case "1011110000" => BCD_output <= "111000010110111101101";
case "1011110001" => BCD_output <= "111000010110111111001";
case "1011110010" => BCD_output <= "111000010110110110011";
case "1011110011" => BCD_output <= "111000010110111011011";
case "1011110100" => BCD_output <= "111000010110111011111";
case "1011110101" => BCD_output <= "111000010110111110000";
case "1011110110" => BCD_output <= "111000010110111111111";
case "1011110111" => BCD_output <= "111000010110111111011";
case "1011111000" => BCD_output <= "111000010111111111110";
case "1011111001" => BCD_output <= "111000010111110110000";
case "1011111010" => BCD_output <= "111000010111111101101";
case "1011111011" => BCD_output <= "111000010111111111001";
case "1011111100" => BCD_output <= "111000010111110110011";
case "1011111101" => BCD_output <= "111000010111111011011";
case "1011111110" => BCD_output <= "111000010111111011111";
case "1011111111" => BCD_output <= "111000010111111110000";
case "1100000000" => BCD_output <= "111000010111111111111";
case "1100000001" => BCD_output <= "111000010111111111011";
case "1100000010" => BCD_output <= "111000011100001111110";
case "1100000011" => BCD_output <= "111000011100000110000";
case "1100000100" => BCD_output <= "111000011100001101101";
case "1100000101" => BCD_output <= "111000011100001111001";
case "1100000110" => BCD_output <= "111000011100000110011";
case "1100000111" => BCD_output <= "111000011100001011011";
case "1100001000" => BCD_output <= "111000011100001011111";
case "1100001001" => BCD_output <= "111000011100001110000";
case "1100001010" => BCD_output <= "111000011100001111111";
case "1100001011" => BCD_output <= "111000011100001111011";
case "1100001100" => BCD_output <= "111000011111111111110";
case "1100001101" => BCD_output <= "111000011111110110000";
case "1100001110" => BCD_output <= "111000011111111101101";
case "1100001111" => BCD_output <= "111000011111111111001";
case "1100010000" => BCD_output <= "111000011111110110011";
case "1100010001" => BCD_output <= "111000011111111011011";
case "1100010010" => BCD_output <= "111000011111111011111";
case "1100010011" => BCD_output <= "111000011111111110000";
case "1100010100" => BCD_output <= "111000011111111111111";
case "1100010101" => BCD_output <= "111000011111111111011";
case "1100010110" => BCD_output <= "111000011110111111110";
case "1100010111" => BCD_output <= "111000011110110110000";
case "1100011000" => BCD_output <= "111000011110111101101";
case "1100011001" => BCD_output <= "111000011110111111001";
case "1100011010" => BCD_output <= "111000011110110110011";
case "1100011011" => BCD_output <= "111000011110111011011";
case "1100011100" => BCD_output <= "111000011110111011111";
case "1100011101" => BCD_output <= "111000011110111110000";
case "1100011110" => BCD_output <= "111000011110111111111";
case "1100011111" => BCD_output <= "111000011110111111011";
case "1100100000" => BCD_output <= "111111111111101111110";
case "1100100001" => BCD_output <= "111111111111100110000";
case "1100100010" => BCD_output <= "111111111111101101101";
case "1100100011" => BCD_output <= "111111111111101111001";
case "1100100100" => BCD_output <= "111111111111100110011";
case "1100100101" => BCD_output <= "111111111111101011011";
case "1100100110" => BCD_output <= "111111111111101011111";
case "1100100111" => BCD_output <= "111111111111101110000";
case "1100101000" => BCD_output <= "111111111111101111111";
case "1100101001" => BCD_output <= "111111111111101111011";
case "1100101010" => BCD_output <= "111111101100001111110";
case "1100101011" => BCD_output <= "111111101100000110000";
case "1100101100" => BCD_output <= "111111101100001101101";
case "1100101101" => BCD_output <= "111111101100001111001";
case "1100101110" => BCD_output <= "111111101100000110011";
case "1100101111" => BCD_output <= "111111101100001011011";
case "1100110000" => BCD_output <= "111111101100001011111";
case "1100110001" => BCD_output <= "111111101100001110000";
case "1100110010" => BCD_output <= "111111101100001111111";
case "1100110011" => BCD_output <= "111111101100001111011";
case "1100110100" => BCD_output <= "111111111011011111110";
case "1100110101" => BCD_output <= "111111111011010110000";
case "1100110110" => BCD_output <= "111111111011011101101";
case "1100110111" => BCD_output <= "111111111011011111001";
case "1100111000" => BCD_output <= "111111111011010110011";
case "1100111001" => BCD_output <= "111111111011011011011";
case "1100111010" => BCD_output <= "111111111011011011111";
case "1100111011" => BCD_output <= "111111111011011110000";
case "1100111100" => BCD_output <= "111111111011011111111";
case "1100111101" => BCD_output <= "111111111011011111011";
case "1100111110" => BCD_output <= "111111111110011111110";
case "1100111111" => BCD_output <= "111111111110010110000";
case "1101000000" => BCD_output <= "111111111110011101101";
case "1101000001" => BCD_output <= "111111111110011111001";
case "1101000010" => BCD_output <= "111111111110010110011";
case "1101000011" => BCD_output <= "111111111110011011011";
case "1101000100" => BCD_output <= "111111111110011011111";
case "1101000101" => BCD_output <= "111111111110011110000";
case "1101000110" => BCD_output <= "111111111110011111111";
case "1101000111" => BCD_output <= "111111111110011111011";
case "1101001000" => BCD_output <= "111111101100111111110";
case "1101001001" => BCD_output <= "111111101100110110000";
case "1101001010" => BCD_output <= "111111101100111101101";
case "1101001011" => BCD_output <= "111111101100111111001";
case "1101001100" => BCD_output <= "111111101100110110011";
case "1101001101" => BCD_output <= "111111101100111011011";
case "1101001110" => BCD_output <= "111111101100111011111";
case "1101001111" => BCD_output <= "111111101100111110000";
case "1101010000" => BCD_output <= "111111101100111111111";
case "1101010001" => BCD_output <= "111111101100111111011";
case "1101010010" => BCD_output <= "111111110110111111110";
case "1101010011" => BCD_output <= "111111110110110110000";
case "1101010100" => BCD_output <= "111111110110111101101";
case "1101010101" => BCD_output <= "111111110110111111001";
case "1101010110" => BCD_output <= "111111110110110110011";
case "1101010111" => BCD_output <= "111111110110111011011";
case "1101011000" => BCD_output <= "111111110110111011111";
case "1101011001" => BCD_output <= "111111110110111110000";
case "1101011010" => BCD_output <= "111111110110111111111";
case "1101011011" => BCD_output <= "111111110110111111011";
case "1101011100" => BCD_output <= "111111110111111111110";
case "1101011101" => BCD_output <= "111111110111110110000";
case "1101011110" => BCD_output <= "111111110111111101101";
case "1101011111" => BCD_output <= "111111110111111111001";
case "1101100000" => BCD_output <= "111111110111110110011";
case "1101100001" => BCD_output <= "111111110111111011011";
case "1101100010" => BCD_output <= "111111110111111011111";
case "1101100011" => BCD_output <= "111111110111111110000";
case "1101100100" => BCD_output <= "111111110111111111111";
case "1101100101" => BCD_output <= "111111110111111111011";
case "1101100110" => BCD_output <= "111111111100001111110";
case "1101100111" => BCD_output <= "111111111100000110000";
case "1101101000" => BCD_output <= "111111111100001101101";
case "1101101001" => BCD_output <= "111111111100001111001";
case "1101101010" => BCD_output <= "111111111100000110011";
case "1101101011" => BCD_output <= "111111111100001011011";
case "1101101100" => BCD_output <= "111111111100001011111";
case "1101101101" => BCD_output <= "111111111100001110000";
case "1101101110" => BCD_output <= "111111111100001111111";
case "1101101111" => BCD_output <= "111111111100001111011";
case "1101110000" => BCD_output <= "111111111111111111110";
case "1101110001" => BCD_output <= "111111111111110110000";
case "1101110010" => BCD_output <= "111111111111111101101";
case "1101110011" => BCD_output <= "111111111111111111001";
case "1101110100" => BCD_output <= "111111111111110110011";
case "1101110101" => BCD_output <= "111111111111111011011";
case "1101110110" => BCD_output <= "111111111111111011111";
case "1101110111" => BCD_output <= "111111111111111110000";
case "1101111000" => BCD_output <= "111111111111111111111";
case "1101111001" => BCD_output <= "111111111111111111011";
case "1101111010" => BCD_output <= "111111111110111111110";
case "1101111011" => BCD_output <= "111111111110110110000";
case "1101111100" => BCD_output <= "111111111110111101101";
case "1101111101" => BCD_output <= "111111111110111111001";
case "1101111110" => BCD_output <= "111111111110110110011";
case "1101111111" => BCD_output <= "111111111110111011011";
case "1110000000" => BCD_output <= "111111111110111011111";
case "1110000001" => BCD_output <= "111111111110111110000";
case "1110000010" => BCD_output <= "111111111110111111111";
case "1110000011" => BCD_output <= "111111111110111111011";
case "1110000100" => BCD_output <= "111101111111101111110";
case "1110000101" => BCD_output <= "111101111111100110000";
case "1110000110" => BCD_output <= "111101111111101101101";
case "1110000111" => BCD_output <= "111101111111101111001";
case "1110001000" => BCD_output <= "111101111111100110011";
case "1110001001" => BCD_output <= "111101111111101011011";
case "1110001010" => BCD_output <= "111101111111101011111";
case "1110001011" => BCD_output <= "111101111111101110000";
case "1110001100" => BCD_output <= "111101111111101111111";
case "1110001101" => BCD_output <= "111101111111101111011";
case "1110001110" => BCD_output <= "111101101100001111110";
case "1110001111" => BCD_output <= "111101101100000110000";
case "1110010000" => BCD_output <= "111101101100001101101";
case "1110010001" => BCD_output <= "111101101100001111001";
case "1110010010" => BCD_output <= "111101101100000110011";
case "1110010011" => BCD_output <= "111101101100001011011";
case "1110010100" => BCD_output <= "111101101100001011111";
case "1110010101" => BCD_output <= "111101101100001110000";
case "1110010110" => BCD_output <= "111101101100001111111";
case "1110010111" => BCD_output <= "111101101100001111011";
case "1110011000" => BCD_output <= "111101111011011111110";
case "1110011001" => BCD_output <= "111101111011010110000";
case "1110011010" => BCD_output <= "111101111011011101101";
case "1110011011" => BCD_output <= "111101111011011111001";
case "1110011100" => BCD_output <= "111101111011010110011";
case "1110011101" => BCD_output <= "111101111011011011011";
case "1110011110" => BCD_output <= "111101111011011011111";
case "1110011111" => BCD_output <= "111101111011011110000";
case "1110100000" => BCD_output <= "111101111011011111111";
case "1110100001" => BCD_output <= "111101111011011111011";
case "1110100010" => BCD_output <= "111101111110011111110";
case "1110100011" => BCD_output <= "111101111110010110000";
case "1110100100" => BCD_output <= "111101111110011101101";
case "1110100101" => BCD_output <= "111101111110011111001";
case "1110100110" => BCD_output <= "111101111110010110011";
case "1110100111" => BCD_output <= "111101111110011011011";
case "1110101000" => BCD_output <= "111101111110011011111";
case "1110101001" => BCD_output <= "111101111110011110000";
case "1110101010" => BCD_output <= "111101111110011111111";
case "1110101011" => BCD_output <= "111101111110011111011";
case "1110101100" => BCD_output <= "111101101100111111110";
case "1110101101" => BCD_output <= "111101101100110110000";
case "1110101110" => BCD_output <= "111101101100111101101";
case "1110101111" => BCD_output <= "111101101100111111001";
case "1110110000" => BCD_output <= "111101101100110110011";
case "1110110001" => BCD_output <= "111101101100111011011";
case "1110110010" => BCD_output <= "111101101100111011111";
case "1110110011" => BCD_output <= "111101101100111110000";
case "1110110100" => BCD_output <= "111101101100111111111";
case "1110110101" => BCD_output <= "111101101100111111011";
case "1110110110" => BCD_output <= "111101110110111111110";
case "1110110111" => BCD_output <= "111101110110110110000";
case "1110111000" => BCD_output <= "111101110110111101101";
case "1110111001" => BCD_output <= "111101110110111111001";
case "1110111010" => BCD_output <= "111101110110110110011";
case "1110111011" => BCD_output <= "111101110110111011011";
case "1110111100" => BCD_output <= "111101110110111011111";
case "1110111101" => BCD_output <= "111101110110111110000";
case "1110111110" => BCD_output <= "111101110110111111111";
case "1110111111" => BCD_output <= "111101110110111111011";
case "1111000000" => BCD_output <= "111101110111111111110";
case "1111000001" => BCD_output <= "111101110111110110000";
case "1111000010" => BCD_output <= "111101110111111101101";
case "1111000011" => BCD_output <= "111101110111111111001";
case "1111000100" => BCD_output <= "111101110111110110011";
case "1111000101" => BCD_output <= "111101110111111011011";
case "1111000110" => BCD_output <= "111101110111111011111";
case "1111000111" => BCD_output <= "111101110111111110000";
case "1111001000" => BCD_output <= "111101110111111111111";
case "1111001001" => BCD_output <= "111101110111111111011";
case "1111001010" => BCD_output <= "111101111100001111110";
case "1111001011" => BCD_output <= "111101111100000110000";
case "1111001100" => BCD_output <= "111101111100001101101";
case "1111001101" => BCD_output <= "111101111100001111001";
case "1111001110" => BCD_output <= "111101111100000110011";
case "1111001111" => BCD_output <= "111101111100001011011";
case "1111010000" => BCD_output <= "111101111100001011111";
case "1111010001" => BCD_output <= "111101111100001110000";
case "1111010010" => BCD_output <= "111101111100001111111";
case "1111010011" => BCD_output <= "111101111100001111011";
case "1111010100" => BCD_output <= "111101111111111111110";
case "1111010101" => BCD_output <= "111101111111110110000";
case "1111010110" => BCD_output <= "111101111111111101101";
case "1111010111" => BCD_output <= "111101111111111111001";
case "1111011000" => BCD_output <= "111101111111110110011";
case "1111011001" => BCD_output <= "111101111111111011011";
case "1111011010" => BCD_output <= "111101111111111011111";
case "1111011011" => BCD_output <= "111101111111111110000";
case "1111011100" => BCD_output <= "111101111111111111111";
case "1111011101" => BCD_output <= "111101111111111111011";
case "1111011110" => BCD_output <= "111101111110111111110";
case "1111011111" => BCD_output <= "111101111110110110000";
case "1111100000" => BCD_output <= "111101111110111101101";
case "1111100001" => BCD_output <= "111101111110111111001";
case "1111100010" => BCD_output <= "111101111110110110011";
case "1111100011" => BCD_output <= "111101111110111011011";
case "1111100100" => BCD_output <= "111101111110111011111";
case "1111100101" => BCD_output <= "111101111110111110000";
case "1111100110" => BCD_output <= "111101111110111111111";
case "1111100111" => BCD_output <= "111101111110111111011";
